// Compatibility wrapper so `` `include "uvm_macros.svh" `` resolves when the
// stub package is used.
`include "uvm_stub_macros.svh"
